// Code your design here
module ternary(input A, input B, output Z);
  assign Z = A > B ? 1 : 0;
endmodule
